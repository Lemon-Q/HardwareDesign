`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/07 13:50:53
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top(
	input wire clk,rst,
	output wire[31:0] writedata,dataadr,
	output wire[3:0] wa
    );

	wire[31:0] pc,instr,readdata;

	mips mips(clk,rst,pc,instr,wa,dataadr,writedata,readdata);
	inst_mem imem(~clk,pc,instr);
	data_mem dmem(~clk,wa,dataadr,writedata,readdata);

endmodule

//git config --global --unset http.proxy